bit [6:0] opcode;
bit branch, mem_read, mem_to_reg, mem_write, alu_src, reg_write;
bit [1:0] alu_op;
