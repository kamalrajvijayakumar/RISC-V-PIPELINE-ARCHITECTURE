logic [4:0]  rdMem;
logic  regWriteMem;
logic [4:0]  rdWb;
logic  regWriteWb;
logic [4:0]  rs1;
logic [4:0]  rs2;
logic [1:0]  ForwardA;
logic [1:0]  ForwardB;
