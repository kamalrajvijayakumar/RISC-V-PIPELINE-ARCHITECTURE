logic clk;
logic reset;
logic [63:0] alu_result;
logic [63:0]adder_ex_out;
logic [63:0]mux_2_out;
logic [4:0]rd;
logic branch_exout;
logic memread_exout;
logic memtoreg_exout;
logic memwrite_exout;
logic regwrite_exout;
logic zero;
       logic [63:0]alu_result_memout;
logic [63:0]adder_ex_out_mem_out;
       logic [63:0] mux_2_out_memout;
       logic [4:0] rd_memout;
logic branch_exout_memout;
logic memread_exout_memout;
logic memtoreg_exout_memout;
logic memwrite_exout_memout;
logic regwrite_exout_memout;
logic zero_memout;