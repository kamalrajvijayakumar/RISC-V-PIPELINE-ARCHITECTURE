bit [63:0] adder_if_out_mux_if_in;
bit [63:0] adder_ex_out_mux_if_in;
bit        and_out;
bit [63:0] mux_if_out_pc_in;
