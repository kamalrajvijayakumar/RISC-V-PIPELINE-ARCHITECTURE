logic [63:0] mux_1_out_alu_in;
logic [63:0] mux_ex_out_alu_in;
logic [3:0]  ALUOp;
logic [63:0] Result;
logic zero;
