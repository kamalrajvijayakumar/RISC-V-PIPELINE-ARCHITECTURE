logic [31:0] instruction_idout;
bit [6:0]  opcode;
bit [4:0]  rd;
bit [2:0]  funct3;
bit [4:0]  rs1;
bit [4:0]  rs2;
bit [6:0]  funct7;
