logic clk;
logic reset;
logic [63:0] pc_out_aim_in;
logic [31:0] instruction;
logic [63:0] pcid_out;
logic [31:0] instruction_idout;