logic clk;
logic reset;
logic [63:0]pcid_out;
logic [63:0]readdata1ex;
logic [63:0]readdata2ex;
logic [63:0] imm_data;
logic [4:0]  rd;
logic [4:0]  rs1;
logic [4:0]  rs2;
logic [31:0] instruction_idout;
logic branch;
logic memread;
logic memtoreg;
logic memwrite;
logic alusrc_in;
logic regwrite;
logic [1:0] aluop_in;
logic [63:0] pcid_exout;
logic [63:0] readdata1ex_out;
logic [63:0] readdata2ex_out;
logic  [63:0] imm_data_exout;
logic [4:0]  rs1_ex;
logic  [4:0]  rs2_ex;
logic [4:0]  rd_ex;
logic [3:0]  instruction_id_exout;
logic branch_exout;
logic memread_exout;
logic memtoreg_exout;
logic memwrite_exout;
logic alusrc;
logic regwrite_exout;
logic [1:0] aluop;
