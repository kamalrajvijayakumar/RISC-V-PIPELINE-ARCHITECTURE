
logic [31:0] alu_out;
logic [31:0] mux3_out_writedata_in;
logic mem_read;
logic mem_write;
logic [31:0] read_data_out_mux5_1_in;
