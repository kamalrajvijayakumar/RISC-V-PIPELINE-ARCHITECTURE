logic [1:0]  ALUOp;
logic [3:0]  func;
logic [3:0]  alu_control;
  