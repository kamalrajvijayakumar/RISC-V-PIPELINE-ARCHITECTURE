logic [63:0] pcid_exout;
logic [63:0] imm_data_exout;
logic [63:0] adder_ex_out_mem_in;
