logic [31:0] instruction_idout;
logic [63:0] imm_data;
