// signals.sv
bit [63:0] pc_out_aim_in;
bit [63:0] adder_if_out_mux_if_in;  
