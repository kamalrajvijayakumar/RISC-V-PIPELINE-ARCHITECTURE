bit clk;
bit reset;
bit [63:0] mux_if_out_pc_in;
bit [63:0] pc_out_aim_in;
