logic branch_exout_memout;
logic zero_memout;
logic and_out;
logic expected;